`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    09:37:30 12/09/2024 
// Design Name: 
// Module Name:    WRITE_MACHINE 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module WRITE_MACHINE(
    input clk,
    input step_en,
    input ack_n,
    output counter_ce,
    output as_n,
    output wr_n,
    output stop_n,
    output in_init,
    output [1:0] wr_state
    );


endmodule
